//-- Alex Grinshpun Apr 2017
//-- Dudy Nov 13 2017
// SystemVerilog version Alex Grinshpun May 2018
// coding convention dudy December 2018
// (c) Technion IIT, Department of Electrical Engineering 2019 


module	background	(	

					input	logic	clk,
					input	logic	resetN,
					input 	logic	[10:0]	pixelX,
					input 	logic	[10:0]	pixelY,

					output	logic	[7:0]	backgroundRGB
);



parameter size = 4;

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 

localparam  int OBJECT_WIDTH_X = 640/size;
localparam  int OBJECT_HEIGHT_Y = 480/size;


logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors = {
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, },
{8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, },
{8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, },
{8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h7B, 8'h9B, 8'h9B, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'hDB, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hBB, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hBB, 8'h9B, 8'hBB, },
{8'hDF, 8'hDB, 8'hBB, 8'hDB, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'hDB, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'hDB, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, },
{8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hFF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDB, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, },
{8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, },
{8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hDE, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hDE, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hDE, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hDF, 8'hDA, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBA, 8'hBE, 8'hBA, 8'hBF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hDF, 8'hDE, 8'hDA, 8'hDA, 8'hDA, 8'hDE, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hDF, 8'hDE, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBA, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hDA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBA, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'h9A, 8'h9A, 8'h9A, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDE, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'h9A, 8'h9A, 8'hBA, 8'hDF, 8'hBA, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hBE, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD8, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'h99, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBF, 8'hDF, 8'hDF, 8'hBA, 8'h99, 8'h9A, 8'h99, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDA, 8'hBA, 8'hBA, 8'hBA, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'h9A, 8'h99, 8'h9A, 8'h9A, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDA, 8'hBA, 8'hBA, 8'hBA, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBE, 8'hDF, 8'hDF, 8'hBA, 8'h99, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDE, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBE, 8'hDF, 8'hDF, 8'h9A, 8'h99, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'h9A, 8'h9A, 8'h9A, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hBE, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBA, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'h9A, 8'h9A, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hBE, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBA, 8'hBA, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hBA, 8'h9A, 8'h9A, 8'hBA, },
{8'h99, 8'h9A, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBE, 8'hBE, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'h99, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'h9A, 8'h99, 8'h99, 8'h96, },
{8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'h9A, 8'h99, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB8, 8'hB8, 8'h98, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h9A, 8'h95, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'h99, 8'h9A, 8'h9A, 8'h95, },
{8'h9A, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBE, 8'hBE, 8'hBA, 8'h9A, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB8, 8'hB8, 8'hB8, 8'h94, 8'hB8, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'h9A, 8'h95, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB8, 8'hB8, 8'hB8, 8'h94, 8'h98, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h96, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'h95, 8'h9A, 8'h9A, 8'h95, },
{8'h95, 8'h9A, 8'h95, 8'h96, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'h9A, 8'h99, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hB8, 8'hB8, 8'hB8, 8'h74, 8'h98, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'h95, 8'h96, 8'h9A, 8'h9A, 8'h9A, 8'h96, 8'h95, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBA, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hB8, 8'hB8, 8'hB8, 8'h94, 8'h94, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h95, 8'h95, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h95, 8'h9A, 8'h95, },
{8'h95, 8'h95, 8'h95, 8'h96, 8'h9A, 8'hBA, 8'hBA, 8'hBA, 8'h9A, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h9A, 8'h9A, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h74, 8'h98, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h9A, 8'h9A, 8'hBA, 8'hBA, 8'h9A, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h9A, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h94, 8'h94, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, },
{8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h96, 8'h95, 8'h99, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h74, 8'h94, 8'hB8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h96, 8'h95, 8'h95, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h74, 8'h94, 8'hB8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, },
{8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h96, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'hB8, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'h99, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h96, 8'h99, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h98, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h96, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, },
{8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hD8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hD8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h99, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h99, 8'hB9, 8'hD9, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hD8, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hD9, 8'hB9, 8'h99, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, },
{8'h99, 8'h99, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hD8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h99, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h98, 8'hB8, 8'hD8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h94, 8'h94, 8'h94, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hD8, 8'hB8, 8'h98, 8'h98, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h98, 8'hB8, 8'hD8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h94, 8'h94, 8'h94, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h94, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h94, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h98, 8'h99, 8'h99, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'h99, 8'h99, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'h74, 8'h94, 8'h94, 8'h94, 8'h94, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, },
{8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, },
{8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, },
{8'h74, 8'h95, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB9, 8'h94, 8'h94, 8'h98, 8'hB8, 8'hD8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB9, 8'h98, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h95, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h99, 8'h74, 8'h94, 8'h99, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB9, 8'hB8, 8'h94, 8'h98, 8'hB8, 8'hD8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB9, 8'hB8, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h95, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h99, 8'h94, 8'h94, 8'h99, 8'h98, },
{8'h95, 8'hB5, 8'h95, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h94, 8'hB4, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h90, 8'h95, 8'hB5, 8'h70, 8'h6C, 8'h70, 8'h70, 8'hB0, 8'h70, 8'h70, 8'h74, 8'h94, 8'hB4, 8'h95, 8'hD9, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'hB4, 8'h94, 8'hD4, 8'hB4, 8'hB5, 8'hB5, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'hB5, 8'hDA, 8'h94, 8'hD4, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h94, 8'h95, 8'h70, 8'h70, 8'h90, 8'hD4, 8'hB5, 8'hDA, 8'h95, 8'hB5, 8'hB5, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'hB4, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h95, 8'hB5, 8'h70, 8'h6C, 8'h70, 8'h70, 8'hB0, 8'h90, 8'h70, 8'h70, 8'h94, 8'hB8, 8'h94, 8'hD9, 8'h95, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'hB4, 8'h94, 8'hB4, 8'hB4, 8'hB5, 8'hB5, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h95, 8'hDA, 8'h95, 8'hB4, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h95, 8'h70, 8'h70, 8'h70, 8'hB4, 8'hB5, 8'hDA, 8'hB5, 8'hB5, 8'hB5, 8'h70, },
{8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h48, 8'h4C, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h44, 8'h44, 8'h44, 8'h48, 8'h48, 8'h4C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h6C, 8'h70, 8'h6C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h4C, 8'h6C, 8'h6C, 8'h70, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h70, 8'h70, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h6C, 8'h6C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h44, 8'h44, 8'h44, 8'h48, 8'h48, 8'h4C, 8'h4C, 8'h6C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h6C, 8'h6C, 8'h70, 8'h4C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h4C, 8'h6C, 8'h4C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h71, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h6C, 8'h6C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h24, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h24, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, }
};

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		backgroundRGB <=	8'hFF;
	end
	else begin
		if ((pixelX  >= 0) &&  (pixelX < 640) && (pixelY  >= 0) &&  (pixelY < 480) )  // inside an external bracket 
			backgroundRGB <= object_colors[pixelY/size][pixelX/size];	//get RGB from the colors table  
		else 
			backgroundRGB <= TRANSPARENT_ENCODING ; // force color to transparent so it will not be displayed 
	end 
end

// decide if to draw the pixel or not 
assign drawingRequest = (backgroundRGB != TRANSPARENT_ENCODING ) ? 1'b0 : 1'b0 ; // get optional transparent command from the bitmpap   


endmodule

