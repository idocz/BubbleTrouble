module background (
    input logic clk,
    input logic resetN,
    input logic [10:0] offsetX, // offset from top left  position 
    input logic [10:0] offsetY,
    input logic InsideRectangle, //input that the pixel is within a bracket 
    output logic drawingRequest, //output that the pixel should be dispalyed 
    output logic [23:0] RGBout //rgb value form the bitmap 
);

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
localparam  int OBJECT_WIDTH_X = 160;
localparam  int OBJECT_HEIGHT_Y = 120;

logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors = {
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, },
{8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, },
{8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, },
{8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, },
{8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h57, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h7B, 8'h9B, 8'h9B, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h77, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, },
{8'hDB, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hBB, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hBB, 8'h9B, 8'hBB, },
{8'hDF, 8'hDB, 8'hBB, 8'hDB, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'hDB, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'hDB, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h9B, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'h9B, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hBB, 8'h9B, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, },
{8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hBB, 8'hBB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hFF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDB, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, },
{8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, },
{8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hDE, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hDE, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hDE, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hDF, 8'hDA, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBA, 8'hBE, 8'hBA, 8'hBF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hDF, 8'hDE, 8'hDA, 8'hDA, 8'hDA, 8'hDE, 8'hDF, 8'hDF, 8'hDB, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hDF, 8'hDE, 8'hDA, 8'hDA, 8'hDA, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBA, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hDA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBA, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDB, 8'h9A, 8'h9A, 8'h9A, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDE, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hDA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'h9A, 8'h9A, 8'hBA, 8'hDF, 8'hBA, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hBE, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD8, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'h99, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hDA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBF, 8'hDF, 8'hDF, 8'hBA, 8'h99, 8'h9A, 8'h99, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDA, 8'hBA, 8'hBA, 8'hBA, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'h9A, 8'h99, 8'h9A, 8'h9A, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDA, 8'hBA, 8'hBA, 8'hBA, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBE, 8'hDF, 8'hDF, 8'hBA, 8'h99, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDF, 8'hDF, 8'hDF, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBA, 8'hBE, 8'hBA, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hDE, 8'hDF, 8'hDF, 8'hDF, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBE, 8'hDF, 8'hDF, 8'h9A, 8'h99, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, 8'hDF, },
{8'h9A, 8'h9A, 8'h9A, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hBE, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBA, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'h9A, 8'h9A, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hBE, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBA, 8'hBA, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hDF, 8'hBA, 8'h9A, 8'h9A, 8'hBA, },
{8'h99, 8'h9A, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBE, 8'hBE, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'h99, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'h9A, 8'h99, 8'h99, 8'h96, },
{8'h9A, 8'h9A, 8'h95, 8'h9A, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'h9A, 8'h99, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hBA, 8'hBA, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB8, 8'hB8, 8'h98, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h9A, 8'h95, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'h99, 8'h9A, 8'h9A, 8'h95, },
{8'h9A, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBE, 8'hBE, 8'hBA, 8'h9A, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB8, 8'hB8, 8'hB8, 8'h94, 8'hB8, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'h9A, 8'h95, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB8, 8'hB8, 8'hB8, 8'h94, 8'h98, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h96, 8'h95, 8'hBA, 8'hBE, 8'hBE, 8'hBA, 8'h95, 8'h9A, 8'h9A, 8'h95, },
{8'h95, 8'h9A, 8'h95, 8'h96, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'h9A, 8'h99, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hB8, 8'hB8, 8'hB8, 8'h74, 8'h98, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'h95, 8'h96, 8'h9A, 8'h9A, 8'h9A, 8'h96, 8'h95, 8'h9A, 8'h95, 8'h96, 8'hBA, 8'hBE, 8'hBE, 8'hBE, 8'hBE, 8'hBA, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hBA, 8'hBE, 8'hBA, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hB8, 8'hB8, 8'hB8, 8'h94, 8'h94, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h95, 8'h95, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h95, 8'h95, 8'h9A, 8'h95, },
{8'h95, 8'h95, 8'h95, 8'h96, 8'h9A, 8'hBA, 8'hBA, 8'hBA, 8'h9A, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h9A, 8'h9A, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h74, 8'h98, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h9A, 8'h9A, 8'hBA, 8'hBA, 8'h9A, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'h9A, 8'h9A, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h94, 8'h94, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, },
{8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h96, 8'h95, 8'h99, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h74, 8'h94, 8'hB8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h96, 8'h95, 8'h95, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h74, 8'h94, 8'hB8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, },
{8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h96, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'hB8, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'h99, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h96, 8'h99, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h98, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h95, 8'h96, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, },
{8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hD8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hD8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'h99, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, 8'h99, 8'hB9, 8'hD9, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hD8, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hD9, 8'hB9, 8'h99, 8'h95, 8'h95, 8'h95, 8'h95, 8'h95, },
{8'h99, 8'h99, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hD8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h99, 8'h99, 8'h99, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h98, 8'hB8, 8'hD8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h94, 8'h94, 8'h94, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hD8, 8'hB8, 8'h98, 8'h98, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h98, 8'hB8, 8'hD8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h94, 8'h94, 8'h94, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hD9, 8'hD9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h94, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h94, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h98, 8'h99, 8'h99, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB9, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'h99, 8'h99, 8'h99, 8'h99, 8'h99, 8'hB9, 8'hB9, 8'hB9, 8'hB9, },
{8'h74, 8'h94, 8'h94, 8'h94, 8'h94, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, },
{8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, },
{8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h98, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, },
{8'h74, 8'h95, 8'h98, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB9, 8'h94, 8'h94, 8'h98, 8'hB8, 8'hD8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB9, 8'h98, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h95, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h94, 8'h99, 8'h74, 8'h94, 8'h99, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'h98, 8'h98, 8'h98, 8'hB8, 8'hB9, 8'hB8, 8'h94, 8'h98, 8'hB8, 8'hD8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'hB8, 8'h98, 8'hB8, 8'hB8, 8'hB8, 8'hB9, 8'hB8, 8'h94, 8'h94, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h95, 8'h94, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'h99, 8'h94, 8'h94, 8'h99, 8'h98, },
{8'h95, 8'hB5, 8'h95, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h94, 8'hB4, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h90, 8'h95, 8'hB5, 8'h70, 8'h6C, 8'h70, 8'h70, 8'hB0, 8'h70, 8'h70, 8'h74, 8'h94, 8'hB4, 8'h95, 8'hD9, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'hB4, 8'h94, 8'hD4, 8'hB4, 8'hB5, 8'hB5, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h94, 8'hB5, 8'hDA, 8'h94, 8'hD4, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h94, 8'h95, 8'h70, 8'h70, 8'h90, 8'hD4, 8'hB5, 8'hDA, 8'h95, 8'hB5, 8'hB5, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'hB4, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h95, 8'hB5, 8'h70, 8'h6C, 8'h70, 8'h70, 8'hB0, 8'h90, 8'h70, 8'h70, 8'h94, 8'hB8, 8'h94, 8'hD9, 8'h95, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'h94, 8'hB4, 8'h94, 8'hB4, 8'hB4, 8'hB5, 8'hB5, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h74, 8'h74, 8'h74, 8'h74, 8'h94, 8'h95, 8'hDA, 8'h95, 8'hB4, 8'h94, 8'h70, 8'h70, 8'h70, 8'h70, 8'h70, 8'h95, 8'h70, 8'h70, 8'h70, 8'hB4, 8'hB5, 8'hDA, 8'hB5, 8'hB5, 8'hB5, 8'h70, },
{8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h48, 8'h4C, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h44, 8'h44, 8'h44, 8'h48, 8'h48, 8'h4C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h6C, 8'h70, 8'h6C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h4C, 8'h6C, 8'h6C, 8'h70, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h70, 8'h70, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h6C, 8'h6C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h44, 8'h44, 8'h44, 8'h48, 8'h48, 8'h4C, 8'h4C, 8'h6C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h6C, 8'h6C, 8'h70, 8'h4C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h48, 8'h4C, 8'h6C, 8'h4C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h71, 8'h4C, 8'h4C, 8'h4C, 8'h6C, 8'h6C, 8'h6C, 8'h6C, 8'h6C, 8'h4C, 8'h4C, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h24, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h24, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h44, 8'h44, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, },
{8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, 8'h24, }
};

wire [7:0] red_sig, green_sig, blue_sig;
assign red_sig     = {object_colors[offsetY][offsetX][7:5] , 5'd0};
assign green_sig   = {object_colors[offsetY][offsetX][4:2] , 5'd0};
assign blue_sig    = {object_colors[offsetY][offsetX][1:0] , 6'd0};


always_ff@(posedge clk)
begin
       RGBout      <= {red_sig,green_sig,blue_sig};
       if (InsideRectangle == 1'b1 ) begin // inside an external bracket 
            if (object_colors[offsetY][offsetX] != TRANSPARENT_ENCODING)
                drawingRequest <= 1'b1;
            else
                drawingRequest <= 1'b0;
       end
       else
            drawingRequest <= 1'b0;
end

endmodule