// (c) Technion IIT, Department of Electrical Engineering 2018 
// Updated by Liat Schwartz March 2019 

// Implements a simple traffic lights controller
// by using state machine with present and next states wvf6

module  presentsController (

	input logic clk, resetN,
	
	input logic dropPresent,
	
	input logic col_player_present1,
	input logic col_rope_present1,
	
	input logic col_player_present2,
	input logic col_rope_present2,
	
	input logic col_player_present3,
	input logic col_rope_present3,
	
	//random present
	input logic [2:0] nxt_present,

	//sec counter
	input logic secClk,
	input logic presentsVisible,
	
	//Visible
	output logic present1Visible,
	output logic present2Visible,
	output logic present3Visible,

	//reset
	output logic present1Reset,
	output logic present2Reset,
	output logic present3Reset,
	
	//presents types
	output logic [1:0] pType1, pType2, pType3,
	
	output logic col_present,
	output logic [1:0] present_type
	
	
);
	
	
enum logic [1:0] {inactive, active} cur_st1, nxt_st1, cur_st2, nxt_st2, cur_st3, nxt_st3;
logic [3:0] timer1, timer2, timer3, nxt_timer1, nxt_timer2, nxt_timer3; 
logic [1:0] nxt_pType1, nxt_pType2, nxt_pType3;
logic nxt_present1Visible, nxt_present2Visible, nxt_present3Visible;
logic nxt_present1Reset, nxt_present2Reset, nxt_present3Reset;
parameter maxTime = 10;


always_ff @(posedge clk or negedge resetN)
begin
   if ( !resetN ) 
	begin // Asynchronic reset	
	
		cur_st1 <= inactive;
		cur_st2 <= inactive;
		cur_st3 <= inactive;
		
		timer1 <= maxTime;
		timer2 <= maxTime;
		timer3 <= maxTime;
		
		pType1 <= 0;
		pType2 <= 0;
		pType3 <= 0;
		
		present1Visible <= 0;
		present2Visible <= 0;
		present3Visible <= 0;

		present1Reset <= 0;
		present2Reset <= 0;
		present3Reset <= 0;
		
	end // asynch
	else
	begin
	
		cur_st1 <= nxt_st1; 
		cur_st2 <= nxt_st2;
		cur_st3 <= nxt_st3;
		
		timer1 <= nxt_timer1;
		timer2 <= nxt_timer2;
		timer3 <= nxt_timer3;
		
		pType1 <= nxt_pType1;
		pType2 <= nxt_pType2;
		pType3 <= nxt_pType3;
		
		present1Visible <= nxt_present1Visible;
		present2Visible <= nxt_present2Visible;
		present3Visible <= nxt_present3Visible;
		
		present1Reset <= nxt_present1Reset;
		present2Reset <= nxt_present2Reset;
		present3Reset <= nxt_present3Reset;
		
	end
end


	
always_comb // Update the next state 1  ////////////////////////////////
begin

		nxt_st1 = cur_st1;	// Set default values
		nxt_st2 = cur_st2;
		nxt_st3 = cur_st3;
		
		nxt_pType1 = pType1;
		nxt_pType2 = pType2;
		nxt_pType3 = pType3;
		
		nxt_timer1 = timer1;
		nxt_timer2 = timer2;
		nxt_timer3 = timer3;
		
		if ( dropPresent == 1'b1 )
		begin
			if (cur_st1 == inactive) begin
				nxt_st1 = active;
				nxt_timer1 = maxTime;
				nxt_pType1 = nxt_present;
			end
				
			else if (cur_st2 == inactive) begin
				nxt_st2 = active;
				nxt_timer2 = maxTime;
				nxt_pType2 = nxt_present;
			end
			
			else if (cur_st3 == inactive) begin
				nxt_st3 = active;
				nxt_timer3 = maxTime;
				nxt_pType3 = nxt_present;
			end
		end

		
		case ( cur_st1 )
		
			active: begin
			
				if ( timer1 > 0 )
				begin
					if ( secClk )
						nxt_timer1 = timer1 - 1;
				end
				else
					nxt_st1 = inactive;
					
				if ( col_rope_present1 || col_player_present1 || presentsVisible == 1'b0 )
					nxt_st1 = inactive;
					
				
			end
		
		endcase
		
		case ( cur_st2 )
		
			active: begin
			
				if ( timer2 > 0 )
				begin
					if ( secClk )
						nxt_timer2 = timer2 - 1;
				end
				else
					nxt_st2 = inactive;
					
				if ( col_rope_present2 || col_player_present2 || presentsVisible == 1'b0 )
					nxt_st2 = inactive;
				
			end
		
		endcase
		
		case ( cur_st3 )
		
			active: begin
			
				if ( timer3 > 0 )
				begin
					if ( secClk )
						nxt_timer3 = timer3 - 1;
				end
				else
					nxt_st3 = inactive;
				
				if ( col_rope_present3 || col_player_present3 || presentsVisible == 1'b0 )
					nxt_st3 = inactive;	
			end
		
		endcase

end // always next state ///////////////////////////////



always_comb // Update the outputs //////////////////////
  begin
  
  	nxt_present1Visible = present1Visible;
	nxt_present2Visible = present2Visible;
	nxt_present3Visible = present3Visible;
	
	nxt_present1Reset = present1Reset;
	nxt_present2Reset = present2Reset;
	nxt_present3Reset = present3Reset;
	
	present_type = 0;
	col_present = 0;
	
	case (cur_st1) // update outputs for present 1
				
		inactive: begin
		
			nxt_present1Visible = 0;
			nxt_present1Reset = 0;
			
		end // inactive
							

		active: begin
		
			nxt_present1Visible = 1;
			nxt_present1Reset = 1;
			
			if ( col_rope_present1 || col_player_present1 )
			begin
					col_present = 1;
					present_type = pType1;
			end
			
		end // active	
	endcase
	
	
	case (cur_st2) // update outputs for present 2
				
		inactive: begin
		
			nxt_present2Visible = 0;
			nxt_present2Reset = 0;
										
		end // inactive
							

		active: begin
		
			nxt_present2Visible = 1;
			nxt_present2Reset = 1;

			if ( col_rope_present2 || col_player_present2 )
			begin
					col_present = 1;
					present_type = pType2;
			end
					
		end // active	
	endcase
	
	case (cur_st3) // update outputs for present3
				
		inactive: begin
		
			nxt_present3Visible = 0;
			nxt_present3Reset = 0;
			
		end // inactive
							

		active: begin
		
			nxt_present3Visible = 1;
			nxt_present3Reset = 1;

			if ( col_rope_present3 || col_player_present3 )
			begin
					col_present = 1;
					present_type = pType3;
			end
					
		end // active	
	endcase
	
end // always outputs //////////////////////////////
	

	
endmodule
