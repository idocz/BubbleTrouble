// (c) Technion IIT, Department of Electrical Engineering 2018 
// Written By Liat Schwartz August 2018 


// Implements the hexadecimal to 7Segment conversion unit
// by using a two-dimensional array

module hexSS
	(
	input logic [3:0] hexin, 		// Data input: hex numbers 0 to f
	input logic darkN, LampTest, 	// Aditional inputs
	output logic [6:0] ss 	// Output for 7Seg display
	);

//Define the transformation table hex to 7Segment	

 
	logic [0:15] [6:0] SevenSeg =	
				'{	7'h40, 
					7'b1111001,
					7'b0100100,
					7'b0110000,
					7'b0011001,
					7'b0010010,
					7'b0000010,
					7'b1111000,
					7'b0000000,
					7'b0011000,
					7'b0001000,
					7'b0000011,
					7'b1000110,
					7'b0100001,
					7'b0000110,
					7'b0001110};
						
 					
	always_comb
	begin
		if (darkN == 1'b0) begin

			ss = 7'b1111111;
		
			end
		else if(LampTest == 1'b1) begin
			ss = SevenSeg[8];
			end
		else begin 
			ss = SevenSeg[hexin];
			end
	end
	

	
endmodule
