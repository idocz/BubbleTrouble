module game (
    input logic clk,
    input logic resetN,
    input logic [10:0] offsetX, // offset from top left  position 
    input logic [10:0] offsetY,
    input logic InsideRectangle, //input that the pixel is within a bracket 
    output logic drawingRequest, //output that the pixel should be dispalyed 
    output logic [23:0] RGBout //rgb value form the bitmap 
);

localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
localparam  int OBJECT_WIDTH_X = 57;
localparam  int OBJECT_HEIGHT_Y = 30;

logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [8-1:0] object_colors = {
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hFF, 8'hFF, 8'hFB, 8'hFB, 8'hFB, 8'hFB, 8'hFF, 8'hFF, 8'hFB, 8'hFB, 8'hFB, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hCD, 8'hCD, 8'hC9, 8'hC9, 8'hED, 8'hE9, 8'hE9, 8'hCD, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hC9, 8'hC9, 8'hC9, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hC9, 8'hC9, 8'hD2, 8'hFF, 8'hCE, 8'hC9, 8'hC9, 8'hC9, 8'hC9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE5, 8'hCD, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hFB, 8'hC9, 8'hE5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA5, 8'hDB, 8'hFF, 8'hFF, 8'hFB, 8'hF6, 8'hC5, 8'hE5, 8'hC5, 8'hC5, 8'hC1, 8'hCE, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hC1, 8'hE5, 8'hC5, 8'hD2, 8'hFB, 8'hFF, 8'hFB, 8'hD6, 8'hC5, 8'hE1, 8'hE1, 8'hCD, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA5, 8'hC5, 8'hC5, 8'hC5, 8'hA9, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hC5, 8'hE5, 8'hC5, 8'hB2, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB2, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hCE, 8'hC5, 8'hE5, 8'hC5, 8'hB2, 8'hCE, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hFF, 8'hFF, 8'hD2, 8'hC5, 8'hE5, 8'hE5, 8'hC5, 8'hCD, 8'hFF, 8'hCD, 8'hC5, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC9, 8'hB6, 8'hD6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hDA, 8'hFF, },
{8'hFF, 8'hFB, 8'hF6, 8'hC9, 8'hE5, 8'hC5, 8'hA5, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hD2, 8'hC9, 8'hE5, 8'hA5, 8'hA9, 8'hFB, 8'hD6, 8'hA5, 8'hC5, 8'hC5, 8'hCE, 8'hFA, 8'hFF, 8'hD2, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hD2, 8'hC9, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hCD, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC5, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, },
{8'hFF, 8'hD6, 8'hE5, 8'hE5, 8'hE5, 8'hB2, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hE5, 8'hE5, 8'hE5, 8'hB2, 8'hDB, 8'hFF, 8'hFF, 8'hDB, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC5, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD6, 8'hFF, 8'hFF, 8'hFB, 8'hCE, 8'hCE, 8'hCE, 8'hCE, 8'hD2, 8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hA9, 8'hC9, 8'hE5, 8'hA9, 8'hAE, 8'hC5, 8'hE5, 8'hE5, 8'hC9, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hED, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hE9, 8'hD2, 8'hFF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD6, 8'hFF, 8'hFF, 8'hD6, 8'hC5, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hDB, 8'hD6, 8'hC5, 8'hB2, 8'hFF, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA9, 8'hDF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hDB, 8'h8E, 8'hC9, 8'hE5, 8'hE5, 8'hC5, 8'hDA, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE9, 8'hE9, 8'hC9, 8'hC9, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hDB, 8'hDB, 8'hB2, 8'hDA, 8'hFB, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC5, 8'hAE, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB6, 8'hFF, },
{8'hFF, 8'hD2, 8'hC5, 8'hC5, 8'hE5, 8'hD2, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hE5, 8'hE5, 8'hC5, 8'hDA, 8'hFA, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC5, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, },
{8'hFF, 8'hFB, 8'hB6, 8'hCD, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hFF, 8'hFF, 8'hD2, 8'hE5, 8'hE5, 8'hC5, 8'hDA, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hAE, 8'hB6, 8'hB6, 8'hB6, 8'hB6, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hD2, 8'hE5, 8'hE5, 8'hC5, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC5, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hA5, 8'hC5, 8'hE5, 8'hD2, 8'hF6, 8'hF6, 8'hCE, 8'hE5, 8'hE5, 8'hC5, 8'hDA, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hEE, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hFF, 8'hED, 8'hE5, 8'hE5, 8'hE5, 8'hCD, 8'hCE, 8'hCE, 8'hEE, 8'hCE, 8'hEE, 8'hF2, 8'hD2, 8'hD6, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hC9, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hF6, 8'hC5, 8'hE5, 8'hC5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hC5, 8'hE5, 8'hC9, 8'hDB, 8'hD2, 8'hC5, 8'hC5, 8'hC5, 8'hDA, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hC9, 8'hC5, 8'hC5, 8'hC9, 8'hFF, 8'hCD, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hA9, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hAD, 8'hAD, 8'hAD, 8'hAD, 8'hAD, 8'hAD, 8'hAD, 8'hAD, 8'hDB, 8'hDB, 8'h8E, 8'h8E, 8'hAE, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hAE, 8'hAE, 8'hB2, 8'hDB, 8'hDB, 8'hB2, 8'hB2, 8'hB2, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hB2, 8'hB2, 8'hB6, 8'hFF, 8'hD6, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hD6, 8'hF2, 8'hF2, 8'hF2, 8'hD2, 8'hD2, 8'hD2, 8'hD2, 8'hD2, 8'hDB, 8'hFF, 8'hFF, 8'hFB, 8'hD2, 8'hCE, 8'hD2, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hCE, 8'hCE, 8'hD2, 8'hFF, 8'hD6, 8'hEE, 8'hEE, 8'hEE, 8'hEE, 8'hEE, 8'hEE, 8'hEE, 8'hEE, 8'hF2, 8'hF2, 8'hF2, 8'hD6, 8'hFF, 8'hD2, 8'hEE, 8'hEE, 8'hF2, 8'hF2, 8'hEE, 8'hF2, 8'hF2, 8'hF2, 8'hF2, 8'hD2, 8'hFF, 8'hFF, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hE5, 8'hE5, 8'hC5, 8'hC5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hCE, 8'hFF, 8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hAD, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hE5, 8'hC5, 8'hD6, 8'hFF, 8'hFF, },
{8'hFF, 8'hF6, 8'hC9, 8'hE9, 8'hE5, 8'hA9, 8'hAE, 8'hAE, 8'h8D, 8'h8D, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hB2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'h8E, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'h92, 8'hB6, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC9, 8'hB2, 8'hB2, 8'hB2, 8'hB2, 8'hAE, 8'hC5, 8'hE5, 8'hC5, 8'hCE, 8'hFF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hE5, 8'hE5, 8'hC9, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hE5, 8'hE5, 8'hCD, 8'hFF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCE, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hE5, 8'hE5, 8'hCD, 8'hFF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hD6, 8'hFF, 8'hD6, 8'hD2, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hD2, 8'hE5, 8'hE5, 8'hE5, 8'hCE, 8'hF2, 8'hD2, 8'hD2, 8'hF2, 8'hEE, 8'hF2, 8'hD2, 8'hD6, 8'hFF, 8'hC9, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hFF, 8'hFF, 8'hD6, 8'hCE, 8'hE5, 8'hE5, 8'hE5, 8'hCD, 8'hFF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hDB, 8'hD2, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hF2, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hC5, 8'hC5, 8'hE5, 8'hC5, 8'hE5, 8'hC5, 8'hA9, 8'hFF, 8'hE9, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hFF, 8'hFF, 8'hC9, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hCD, 8'hFF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hFB, 8'hAD, 8'hC9, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hE9, 8'hE5, 8'hE5, 8'hE5, 8'hAD, 8'hB2, 8'hDF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hAD, 8'hB2, 8'hAE, 8'hAE, 8'hAE, 8'hAE, 8'hAE, 8'hAE, 8'hB2, 8'hFF, 8'hE9, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hED, 8'hCD, 8'hE5, 8'hE5, 8'hA9, 8'hAE, 8'hAE, 8'hB2, 8'hFF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hE5, 8'hE5, 8'hE5, 8'hD6, 8'hFF, 8'hFF, 8'hD2, 8'hC5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hA5, 8'hD6, 8'hFF, 8'hFF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hD2, 8'hFB, 8'hFF, 8'hFF, 8'hFF, },
{8'hFF, 8'hF6, 8'hE5, 8'hE5, 8'hE5, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hE5, 8'hE5, 8'hE5, 8'hD6, 8'hFF, 8'hFF, 8'hDB, 8'hB2, 8'hC9, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hCD, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hF2, 8'hE5, 8'hE5, 8'hC5, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hE9, 8'hE5, 8'hE5, 8'hC9, 8'hB6, 8'hCD, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hFF, 8'hFF, },
{8'hFF, 8'hD6, 8'hC5, 8'hC5, 8'hE5, 8'hCE, 8'hFB, 8'hFA, 8'hFB, 8'hFB, 8'hEE, 8'hE5, 8'hC5, 8'hA9, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hCD, 8'hA5, 8'hE5, 8'hC5, 8'hA9, 8'hB2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hF2, 8'hE5, 8'hE5, 8'hE5, 8'hCE, 8'hF6, 8'hF2, 8'hF6, 8'hF6, 8'hF6, 8'hF2, 8'hF2, 8'hFB, 8'hFF, 8'hE9, 8'hE5, 8'hE5, 8'hC9, 8'hFF, 8'hD6, 8'hA9, 8'hE5, 8'hE5, 8'hE5, 8'hC5, 8'hD2, 8'hFB, 8'hFF, },
{8'hFF, 8'hFF, 8'hB6, 8'hCD, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hAE, 8'hB6, 8'hDB, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hD6, 8'hC5, 8'hC9, 8'hDB, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hC5, 8'hE5, 8'hC9, 8'hFF, 8'hCD, 8'hE5, 8'hE5, 8'hC9, 8'hDB, 8'hFF, 8'hDB, 8'hCD, 8'hE5, 8'hE5, 8'hE5, 8'hE5, 8'hC9, 8'hDF, },
{8'hFF, 8'hFF, 8'hFF, 8'hD2, 8'hA9, 8'hA9, 8'hA9, 8'hA9, 8'hA9, 8'hA9, 8'hA9, 8'hA9, 8'hD6, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hAD, 8'h8E, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDA, 8'h8E, 8'h8E, 8'h8E, 8'h8E, 8'h8E, 8'h8D, 8'h8D, 8'h8D, 8'h8D, 8'hAE, 8'h8D, 8'hB2, 8'hFF, 8'hD6, 8'h8D, 8'h8D, 8'h8E, 8'hDB, 8'hFF, 8'hFF, 8'hD6, 8'hAD, 8'h8D, 8'h8D, 8'h89, 8'hAE, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDB, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hDF, 8'hDF, 8'hDF, 8'hFF, 8'hFF, },
{8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, }
};

wire [7:0] red_sig, green_sig, blue_sig;
assign red_sig     = {object_colors[offsetY][offsetX][7:5] , 5'd0};
assign green_sig   = {object_colors[offsetY][offsetX][4:2] , 5'd0};
assign blue_sig    = {object_colors[offsetY][offsetX][1:0] , 6'd0};


always_ff@(posedge clk)
begin
       RGBout      <= {red_sig,green_sig,blue_sig};
       if (InsideRectangle == 1'b1 ) begin // inside an external bracket 
            if (object_colors[offsetY][offsetX] != TRANSPARENT_ENCODING)
                drawingRequest <= 1'b1;
            else
                drawingRequest <= 1'b0;
       end
       else
            drawingRequest <= 1'b0;
end

endmodule